module or2 (
    input wire a,  // Input A
    input wire b,  // Input B
    output wire y  // Output Y
);

    assign y = a | b;  // Bitwise OR operation

endmodule
