module buff (
    input wire I,  // Input A
    output wire Z  // Output Y
);

    assign Z = I;  // Directly connect input to output

endmodule
